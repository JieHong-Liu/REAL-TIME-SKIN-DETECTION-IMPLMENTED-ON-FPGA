module secondScan();
endmodule	